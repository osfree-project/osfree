# edlin.sv - Swedish-language messages file
#
# Author: Gregory Pietsch
#
# DESCRIPTION:
#
# This file contains #defines for all the message strings in edlin.
# For internationalization fun, just translate the messages in this
# file.
# Swedish translation Oct 2006 /A.J

1.0:Jj
1.1:: \b
1.2:OK? \b
1.3:Input Error
1.4:%s: %lu rad inl�st\n
1.5:%s: %lu rader inl�sta\n
1.6:%s: %lu rad skriven\n
1.7:%s: %lu rader skrivna\n
1.8:%lu:%c%s\n
1.9:Tryck <enter> 
1.10:%lu: \b
1.11:hittades ej
1.12:%lu: %s\n
1.13:\nedlin har f�ljande (engelska) kommandon:\n
1.14:#                 editera en rad        [#],[#],#m        move
1.15:a                 append                [#][,#]p          page
1.16:[#],[#],#,[#]c    copy                  q                 quit
1.17:[#][,#]d          delete                [#][,#][?]r$,$    replace
1.18:e<>               end (write & quit)    [#][,#][?]s$      s�k
1.19:[#]i              insert                [#]t<>            transfer
1.20:[#][,#]l          lista                 [#]w<>            write\n
1.21:d�r $ �r en str�ng, <> �r ett filnamn,
1.22:# �r ett radnummer (.=aktuell rad, $=sista raden,
1.23: uttryck med +/- kan anv�ndas)\n
1.24:, copyright (c) 2003 Gregory Pietsch
1.25:This program comes with ABSOLUTELY NO WARRANTY.
1.26:It is free software, and you are welcome to redistribute it
1.27:under the terms of the GNU General Public License -- either
1.28:version 2 of the license, or, at your option, any later
1.29:version.\n
1.30:Slut p� minne
1.31:Felaktig Str�ngl�ngd
1.32:Felaktig Str�ngposition
1.33:F�rst�r ej, skriv ? f�r hj�lp.
1.34:Filnamn saknas
1.35:F�r stor buffert
1.36:Ogiltig buffertposition
1.37:ERROR: %s\n

# END OF FILE
